magic
tech sky130A
timestamp 1737732226
<< locali >>
rect -956 -202 -860 -102
rect -380 -202 -284 -110
rect -998 -205 -284 -202
rect -998 -295 -761 -205
rect -671 -295 -284 -205
rect -998 -298 -284 -295
<< viali >>
rect -761 -295 -671 -205
<< metal1 >>
rect -828 916 -796 1466
rect -828 -166 -796 884
rect -764 -205 -668 1698
rect -548 1652 -252 1748
rect -348 1248 -252 1652
rect -548 1152 -252 1248
rect -566 916 -534 919
rect -566 881 -534 884
rect -348 548 -252 1152
rect -572 452 -252 548
rect -348 194 -252 452
rect -572 98 -252 194
rect -764 -295 -761 -205
rect -671 -295 -668 -205
rect -764 -301 -668 -295
<< via1 >>
rect -828 884 -796 916
rect -566 884 -534 916
<< metal2 >>
rect -1066 884 -828 916
rect -796 884 -566 916
rect -534 884 -531 916
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1737728888
transform 1 0 -908 0 1 1414
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1737728888
transform 1 0 -908 0 1 -186
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1737728888
transform 1 0 -908 0 1 214
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1737728888
transform 1 0 -908 0 1 1014
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1737728888
transform 1 0 -908 0 1 614
box -92 -64 668 464
<< labels >>
flabel locali -998 -298 -902 -202 0 FreeSans 800 0 0 0 VSS
port 0 nsew
flabel metal2 -1066 884 -1034 916 0 FreeSans 800 0 0 0 IBPS_5U
port 1 nsew
flabel metal1 -348 98 -252 1748 0 FreeSans 800 0 0 0 IBNS_20U
port 3 nsew
<< end >>
